`ifndef PARAMS_VH
`define PARAMS_VH

`define  FPU_OP_ADD   6'b000_001   
`define  FPU_OP_SUB   6'b000_010   
`define  FPU_OP_MULT  6'b000_011    
`define size_Fp_fmt 3

`endif