module top_core_swc_wrapper (
    input wire hclk,
    input wire hrstn,
    input wire itcm_hready,
    input wire itcm_hresp,
    input wire [31:0] itcm_hrdata,
    input wire itcm_ready,
    input wire dtcm_hready,
    input wire dtcm_hresp,
    input wire [31:0] dtcm_hrdata,
    input wire [3:0] cycle_cnt,
    output wire ifu_dec_stall,
    output wire pc_write,
    output wire [31:0] pc_wdata,
    output wire dec_or,
    output wire [4:0] exu_load_rd,
    output wire [31:0] exu_load_base_addr,
    output wire [31:0] exu_load_offset,
    output wire exu_load_sext,
    output wire [1:0] exu_load_size,
    output wire exu_load_en,
    output wire [31:0] exu_store_addr,
    output wire [31:0] exu_store_data,
    output wire [1:0] exu_store_size,
    output wire exu_store_en,
    output wire [4:0] reg_waddr,
    output wire [31:0] reg_wdata,
    output wire reg_wen,
    output wire [4:0] reg_raddr_1,
    output wire [31:0] reg_rdata_1,
    output wire reg_ren_1,
    output wire [4:0] reg_raddr_2,
    output wire [31:0] reg_rdata_2,
    output wire reg_ren_2,
    output wire pc_write_out,
    output wire [31:0] pc_wdata_out,
    output wire [31:0] mau_haddr,
    output wire mau_hwrite,
    output wire [31:0] mau_hwdata,
    output wire [2:0] mau_hsize,
    output wire [2:0] mau_hburst,
    output wire [6:0] mau_hprot,
    output wire [1:0] mau_htrans,
    output wire mau_hmastlock,
    output wire [4:0] mau_load_rd,
    output wire [31:0] mau_load_data,
    output wire mau_load_en,
    output wire [31:0] ifu_haddr,
    output wire [31:0] ifu_hwdata,
    output wire [31:0] ifu_pc,
    output wire [31:0] ifu_inst_out,
    output wire dec_add,
    output wire [31:0] dec_inst_out,
    output wire [4:0] dec_rs1,
    output wire [4:0] dec_rs2,
    output wire [4:0] dec_rd,
    output wire dec_lw,
    output wire [31:0] regfile [31:0]
);

    top_core_swc dut (
        .hclk(hclk),
        .hrstn(hrstn),
        .itcm_hready(itcm_hready),
        .itcm_hresp(itcm_hresp),
        .itcm_hrdata(itcm_hrdata),
        .itcm_ready(itcm_ready),
        .dtcm_hready(dtcm_hready),
        .dtcm_hresp(dtcm_hresp),
        .dtcm_hrdata(dtcm_hrdata),
        .cycle_cnt(cycle_cnt),
        .ifu_dec_stall(ifu_dec_stall),
        .pc_write(pc_write),
        .pc_wdata(pc_wdata),
        .dec_or(dec_or),
        .exu_load_rd(exu_load_rd),
        .exu_load_base_addr(exu_load_base_addr),
        .exu_load_offset(exu_load_offset),
        .exu_load_sext(exu_load_sext),
        .exu_load_size(exu_load_size),
        .exu_load_en(exu_load_en),
        .exu_store_addr(exu_store_addr),
        .exu_store_data(exu_store_data),
        .exu_store_size(exu_store_size),
        .exu_store_en(exu_store_en),
        .reg_waddr(reg_waddr),
        .reg_wdata(reg_wdata),
        .reg_wen(reg_wen),
        .reg_raddr_1(reg_raddr_1),
        .reg_rdata_1(reg_rdata_1),
        .reg_ren_1(reg_ren_1),
        .reg_raddr_2(reg_raddr_2),
        .reg_rdata_2(reg_rdata_2),
        .reg_ren_2(reg_ren_2),
        .pc_write_out(pc_write_out),
        .pc_wdata_out(pc_wdata_out),
        .mau_haddr(mau_haddr),
        .mau_hwrite(mau_hwrite),
        .mau_hwdata(mau_hwdata),
        .mau_hsize(mau_hsize),
        .mau_hburst(mau_hburst),
        .mau_hprot(mau_hprot),
        .mau_htrans(mau_htrans),
        .mau_hmastlock(mau_hmastlock),
        .mau_load_rd(mau_load_rd),
        .mau_load_data(mau_load_data),
        .mau_load_en(mau_load_en),
        .ifu_haddr(ifu_haddr),
        .ifu_hwdata(ifu_hwdata),
        .ifu_pc(ifu_pc),
        .ifu_inst_out(ifu_inst_out),
        .dec_add(dec_add),
        .dec_inst_out(dec_inst_out),
        .dec_rs1(dec_rs1),
        .dec_rs2(dec_rs2),
        .dec_rd(dec_rd),
        .dec_lw(dec_lw),
        .[31:0]([31:0])
    );
    initial begin
        $dumpfile("./vcds/top_core_swc.vcd");
        $dumpvars(0, top_core_swc_wrapper);
    end
endmodule
